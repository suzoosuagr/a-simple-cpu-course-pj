// Core
// Top-level

module core(clk, CLB);
input wire clk, CLB;

wire 